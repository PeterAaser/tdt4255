library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use work.Defs.ALL;

entity IDEX is
    Generic(
        DATA_WIDTH : integer := 32
    );
    Port ( clk                  : in STD_LOGIC;
           stall                : in STD_LOGIC;
           ControlSignals_in    : in control_signals_t;
           ReadData1_in         : in STD_LOGIC_VECTOR(DATA_WIDTH-1 downto 0);
           ReadData2_in         : in STD_LOGIC_VECTOR(DATA_WIDTH-1 downto 0);
           Immidiate_in         : in immediate_t;
           RegT_in              : in reg_t;
           RegD_in              : in reg_t;
           ControlSignals_out   : out control_signals_t;
           ReadData1_out        : out STD_LOGIC_VECTOR(DATA_WIDTH-1 downto 0);
           ReadData2_out        : out STD_LOGIC_VECTOR(DATA_WIDTH-1 downto 0);
           Immidiate_out        : out STD_LOGIC_VECTOR(DATA_WIDTH-1 downto 0);
           Reg_out             : out reg_t
   );
end IDEX;

architecture Behavioral of IDEX is
begin
    propagate : process(clk)
    begin
        if (rising_edge(clk) and stall = '0')then
           ControlSignals_out <= ControlSignals_in;
           ReadData1_out <= ReadData1_in;
           ReadData2_out <= ReadData2_in;
           Immidiate_out <= std_logic_vector(resize(signed(Immidiate_in), 32));
           if (ControlSignals_in.RegDst = REGT) then
                Reg_out <= RegT_in;
           else
                Reg_out <= RegD_in;
           end if;
       end if;
    end process;
end Behavioral;

