
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all

entity Hazard_detection is

end Hazard_detection;

architecture Behavioral of Hazard_detection is

begin


end Behavioral;

