library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;
use work.defs.all;


entity InstructionDecoder is
end InstructionDecoder;

architecture Behavioral of InstructionDecoder is

begin


end Behavioral;

